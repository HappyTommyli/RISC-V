module csr_reg (
    input wire         clk,          // Clock signal 
    input wire         rst,          // Asynchronous reset 
    input wire [11:0]  csr_addr,     // 12-bit CSR address 
    input wire         csr_write_enable, // Write enable 
    input wire [1:0]   csr_op,       // Operation type (00=CSRRW, 01=CSRRS, 10=CSRRC, 11=immediate variants)
    input wire [2:0]   csr_funct3,   // funct3 field from instruction 
    input wire [31:0]  rs1_data,     // rs1 register data 
    input wire [4:0]   csr_imm,      // 5-bit immediate 
    output reg [31:0]  csr_rdata     // Read CSR value 
);
reg [31:0] mstatus;  // Machine Status Register 
reg [31:0] mie;      // Machine Interrupt Enable Register 
reg [31:0] mtvec;    // Machine Trap Vector Register 
wire [31:0] imm_extended = {27'b0, csr_imm};
always @(*) begin
    case (csr_addr)
        12'h300: csr_rdata = mstatus;
        12'h304: csr_rdata = mie;
        12'h305: csr_rdata = mtvec;
        default: csr_rdata = 32'h0;  // Unimplemented CSRs return 0
    endcase
end
always @(posedge clk or posedge rst) begin
    if (rst) begin
        // Reset to RISC-V default values
        mstatus <= 32'h0;
        mie     <= 32'h0;
        mtvec   <= 32'h0;
    end else if (csr_write_enable) begin
        case (csr_addr)
            12'h300: begin  
                case (csr_op)
                    2'b00: mstatus <= rs1_data;                  // CSRRW
                    2'b01: mstatus <= mstatus | rs1_data;        // CSRRS
                    2'b10: mstatus <= mstatus & (~rs1_data);     // CSRRC
                    2'b11: begin  
                        case (csr_funct3)
                            3'b101: mstatus <= imm_extended;     // CSRRWI
                            3'b110: mstatus <= mstatus | imm_extended;  // CSRRSI
                            3'b111: mstatus <= mstatus & (~imm_extended); // CSRRCI
                            default: ;  // no operation
                        endcase
                    end
                endcase
            end

            12'h304: begin  
                case (csr_op)
                    2'b00: mie <= rs1_data;                      // CSRRW
                    2'b01: mie <= mie | rs1_data;                // CSRRS
                    2'b10: mie <= mie & (~rs1_data);             // CSRRC
                    2'b11: begin  // Immediate variants
                        case (csr_funct3)
                            3'b101: mie <= imm_extended;         // CSRRWI
                            3'b110: mie <= mie | imm_extended;    // CSRRSI
                            3'b111: mie <= mie & (~imm_extended); // CSRRCI
                            default: ;
                        endcase
                    end
                endcase
            end

            12'h305: begin  
                case (csr_op)
                    2'b00: mtvec <= rs1_data;                    // CSRRW
                    2'b01: mtvec <= mtvec | rs1_data;            // CSRRS
                    2'b10: mtvec <= mtvec & (~rs1_data);         // CSRRC
                    2'b11: begin  // Immediate variants
                        case (csr_funct3)
                            3'b101: mtvec <= imm_extended;       // CSRRWI
                            3'b110: mtvec <= mtvec | imm_extended;  // CSRRSI
                            3'b111: mtvec <= mtvec & (~imm_extended); // CSRRCI
                            default: ;
                        endcase
                    end
                endcase
            end

            default: ;  
        endcase
    end
end

endmodule