module control_unit ( 
    input wire [31:0] instruction, 
    output reg reg_write, 
    output reg mem_to_reg, 
    output reg mem_write, 
    output reg mem_read, 
    output reg alu_src, 
    output reg alu_src1,
    output reg [3:0] alu_op, 
    output reg branch, 
    output reg jump, 
    output reg jalr_enable, 
    output reg [11:0] csr_addr, 
    output reg csr_write_enable, 
    output reg [1:0] csr_op, 
    output reg [4:0] csr_imm, 
    output reg [2:0] csr_funct3 
);
    wire [6:0] opcode = instruction[6:0];
    wire [2:0] funct3 = instruction[14:12];
    wire [6:0] funct7 = instruction[31:25];
    wire [11:0] csr_addr_raw = instruction[31:20];
    wire [4:0] csr_imm_raw = instruction[19:15];

    always @(*) begin
        // Defaults
        reg_write = 0; mem_to_reg = 0; mem_write = 0; mem_read = 0;
        alu_src = 0; alu_src1 = 0; alu_op = 4'b0000;
        branch = 0; jump = 0; jalr_enable = 0;
        csr_addr = 0; csr_write_enable = 0; csr_op = 0; csr_imm = 0; csr_funct3 = 0;

        case (opcode)
            7'b0110011: begin // R-type
                reg_write = 1; alu_src = 0;
                case ({funct7, funct3})
                    10'b0000000000: alu_op = 4'b0000; // ADD
                    10'b0100000000: alu_op = 4'b0001; // SUB
                    10'b0000000001: alu_op = 4'b0100; // SLL
                    10'b0000000010: alu_op = 4'b0010; // SLT
                    10'b0000000011: alu_op = 4'b0011; // SLTU
                    10'b0000000100: alu_op = 4'b0101; // XOR
                    10'b0000000101: alu_op = 4'b0110; // SRL
                    10'b0100000101: alu_op = 4'b0111; // SRA
                    10'b0000000110: alu_op = 4'b1000; // OR
                    10'b0000000111: alu_op = 4'b1001; // AND
                    default: alu_op = 4'b1111;
                endcase
            end
            7'b0010011: begin // I-type Arithmetic
                reg_write = 1; alu_src = 1;
                case (funct3)
                    3'b000: alu_op = 4'b0000; // ADDI
                    3'b001: alu_op = 4'b0100; // SLLI
                    3'b010: alu_op = 4'b0010; // SLTI
                    3'b011: alu_op = 4'b0011; // SLTIU
                    3'b100: alu_op = 4'b0101; // XORI
                    3'b101: alu_op = (funct7 == 7'b0100000) ? 4'b0111 : 4'b0110; // SRAI or SRLI
                    3'b110: alu_op = 4'b1000; // ORI
                    3'b111: alu_op = 4'b1001; // ANDI
                    default: alu_op = 4'b1111;
                endcase
            end
            7'b0000011: begin // Loads
                reg_write = 1; mem_to_reg = 1; mem_read = 1; alu_src = 1;
                alu_op = 4'b0000; // ADD
            end
            7'b0100011: begin // Stores
                mem_write = 1; alu_src = 1;
                alu_op = 4'b0000; // ADD
            end
            7'b1100011: begin // Branches
                branch = 1;
                case (funct3)
                    3'b000: alu_op = 4'b0001; // BEQ (use SUB)
                    3'b001: alu_op = 4'b0001; // BNE (use SUB)
                    3'b100: alu_op = 4'b0010; // BLT (use SLT)
                    3'b101: alu_op = 4'b1011; // BGE (use logic >=)
                    3'b110: alu_op = 4'b0011; // BLTU (use SLTU)
                    3'b111: alu_op = 4'b0011; // BGEU (use SLTU logic, inverted in PC_update)
                    default: alu_op = 4'b1111;
                endcase
            end
            7'b1101111: begin // JAL
                reg_write = 1; jump = 1; alu_op = 4'b1010;
            end
            7'b1100111: begin // JALR
                reg_write = 1; jump = 1; jalr_enable = 1; alu_src = 1; alu_op = 4'b0000; // ADD
            end
            7'b0110111: begin // LUI
                reg_write = 1; alu_src = 1; alu_src1 = 0; alu_op = 4'b0000; // ADD (rs1 forced to 0 in EX)
            end
            7'b0010111: begin // AUIPC
                reg_write = 1; alu_src = 1; alu_src1 = 1; alu_op = 4'b0000; // ADD (PC + imm)
            end
            default: alu_op = 4'b1111;
        endcase
    end
endmodule
