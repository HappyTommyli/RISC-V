module PC_update (
    input [31:0] rs1_data, input jump;input branch, input [31:0]pc_address,input [31:0]imm,input zero,output reg next_pc
  );



endmodule
